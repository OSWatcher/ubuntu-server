{
  "MIME": "text/plain",
  "inode_type": "REG",
  "magic_type": "ASCII text",
  "mode": "-rw-r--r--",
  "sha1": "a66dec61fb40335751ea3833a4e4a7c87c97919a"
}