{
  "MIME": "text/plain",
  "inode_type": "REG",
  "magic_type": "UTF-8 Unicode text, with very long lines",
  "mode": "-rw-r--r--",
  "sha1": "545398edfe38a0ce1df93cad88daff74d7efcfe6"
}